bind arbiter check_arbiter arbiter_inst(.*);
